module matrix_operaRTL_1cycle
#(
  parameter number = 9
  )
(
  input
  input   logic   [31:0]  Ix    [number-1:0],
  input   logic   [31:0]  Iy    [number-1:0],
  input   logic   [31:0]  It    [number-1:0],


  );
